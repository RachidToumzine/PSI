--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   18:35:40 05/31/2019
-- Design Name:   
-- Module Name:   /home/toumzine/Bureau/WORK/toumzinecompilateur/process/shema_general_test.vhd
-- Project Name:  process
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: shema_generale
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY shema_general_test IS
END shema_general_test;
 
ARCHITECTURE behavior OF shema_general_test IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT shema_generale
    PORT(
         clk : IN  std_logic;
         rst : IN  std_logic;
         dec_signal : IN  std_logic_vector(31 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal clk : std_logic := '0';
   signal rst : std_logic := '0';
   signal dec_signal : std_logic_vector(31 downto 0) := (others => '0');

   -- Clock period definitions
   constant clk_period : time := 100 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: shema_generale PORT MAP (
          clk => clk,
          rst => rst,
          dec_signal => dec_signal
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	
		
		dec_signal <= x"0601ABCD";
      wait for clk_period;
		
		dec_signal <= x"06020001";
      wait for clk_period;
		
		dec_signal <= x"00000000";
		wait for clk_period*5;
		
		dec_signal <= x"05060100";
		wait for clk_period;

		dec_signal <= x"01010102";
		wait for clk_period*5;

      -- insert stimulus here 

      wait;
		
		-------
		
				
	
	--------------
   end process;

END;
